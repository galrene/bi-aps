module testbench();
	reg         clk;
	reg         reset;
	wire [31:0] data_to_mem, address_to_mem;
	wire        write_enable;

	top simulated_system (clk, reset, data_to_mem, address_to_mem, write_enable);

	initial	begin
		$dumpfile("test.out");
		$dumpvars;
		reset<=1; # 2; reset<=0;
		$writememh ("memfile_data_after_simulation.hex",simulated_system.dmem.RAM,0,63);
		#100;
		$finish;
	end

	// generate clock
	always	begin
		clk<=1; # 1; clk<=0; # 1;
	end
endmodule